magic
tech sky130B
magscale 1 2
timestamp 1733623679
<< pwell >>
rect -296 -279 296 279
<< nmos >>
rect -100 -131 100 69
<< ndiff >>
rect -158 57 -100 69
rect -158 -119 -146 57
rect -112 -119 -100 57
rect -158 -131 -100 -119
rect 100 57 158 69
rect 100 -119 112 57
rect 146 -119 158 57
rect 100 -131 158 -119
<< ndiffc >>
rect -146 -119 -112 57
rect 112 -119 146 57
<< psubdiff >>
rect -260 209 260 243
rect -260 -209 -226 209
rect 226 -209 260 209
rect -260 -243 -164 -209
rect 164 -243 260 -209
<< psubdiffcont >>
rect -164 -243 164 -209
<< poly >>
rect -100 141 100 157
rect -100 107 -84 141
rect 84 107 100 141
rect -100 69 100 107
rect -100 -157 100 -131
<< polycont >>
rect -84 107 84 141
<< locali >>
rect -100 107 -84 141
rect 84 107 100 141
rect -146 57 -112 73
rect -146 -135 -112 -119
rect 112 57 146 73
rect 112 -135 146 -119
rect -180 -243 -164 -209
rect 164 -243 180 -209
<< viali >>
rect -84 107 84 141
rect -146 -119 -112 57
rect 112 -84 146 22
<< metal1 >>
rect -96 141 96 147
rect -96 107 -84 141
rect 84 107 96 141
rect -96 101 96 107
rect -152 57 -106 69
rect -152 -119 -146 57
rect -112 -119 -106 57
rect 106 22 152 34
rect 106 -84 112 22
rect 146 -84 152 22
rect 106 -96 152 -84
rect -152 -131 -106 -119
<< labels >>
flabel metal1 s -2 128 -2 128 0 FreeSans 320 0 0 0 G
port 0 nsew
flabel metal1 s -128 -40 -128 -40 0 FreeSans 320 0 0 0 D
port 1 nsew
flabel metal1 s 128 -38 128 -38 0 FreeSans 320 0 0 0 S
port 2 nsew
flabel locali s 2 -226 2 -226 0 FreeSans 320 0 0 0 B
port 4 nsew
<< properties >>
string FIXED_BBOX -243 -226 243 226
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 1 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 0 gbc 1 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 0 viasrc 60 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
