magic
tech sky130B
magscale 1 2
timestamp 1733616804
<< nwell >>
rect -211 -334 211 334
<< pmos >>
rect -15 -186 15 114
<< pdiff >>
rect -73 102 -15 114
rect -73 -174 -61 102
rect -27 -174 -15 102
rect -73 -186 -15 -174
rect 15 102 73 114
rect 15 -174 27 102
rect 61 -174 73 102
rect 15 -186 73 -174
<< pdiffc >>
rect -61 -174 -27 102
rect 27 -174 61 102
<< nsubdiff >>
rect -175 264 -79 298
rect 79 264 175 298
rect -175 -264 -141 264
rect 141 -264 175 264
rect -175 -298 175 -264
<< nsubdiffcont >>
rect -79 264 79 298
<< poly >>
rect -33 195 33 211
rect -33 161 -17 195
rect 17 161 33 195
rect -33 145 33 161
rect -15 114 15 145
rect -15 -212 15 -186
<< polycont >>
rect -17 161 17 195
<< locali >>
rect -95 264 -79 298
rect 79 264 95 298
rect -33 161 -17 195
rect 17 161 33 195
rect -61 102 -27 118
rect -61 -190 -27 -174
rect 27 102 61 118
rect 27 -190 61 -174
<< viali >>
rect -17 161 17 195
rect -61 -174 -27 102
rect 27 -119 61 47
<< metal1 >>
rect -32 195 36 208
rect -32 161 -17 195
rect 17 161 36 195
rect -32 146 36 161
rect -67 102 -21 114
rect -67 -174 -61 102
rect -27 -174 -21 102
rect 21 47 67 59
rect 21 -119 27 47
rect 61 -119 67 47
rect 21 -131 67 -119
rect -67 -186 -21 -174
<< labels >>
flabel metal1 s 2 178 2 178 0 FreeSans 320 0 0 0 G
port 0 nsew
flabel metal1 s -44 -34 -44 -34 0 FreeSans 320 0 0 0 D
port 1 nsew
flabel metal1 s 44 -40 44 -40 0 FreeSans 320 0 0 0 S
port 2 nsew
flabel locali s 0 280 0 280 0 FreeSans 320 0 0 0 B
port 4 nsew
<< properties >>
string FIXED_BBOX -158 -281 158 281
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.5 l 0.15 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 0 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 60 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
