magic
tech sky130B
magscale 1 2
timestamp 1733623679
use sky130_fd_pr__nfet_01v8_H4FFAF  sky130_fd_pr__nfet_01v8_H4FFAF_0
timestamp 1733623679
transform 1 0 243 0 1 226
box -296 -279 296 279
<< end >>
