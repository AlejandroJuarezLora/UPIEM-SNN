magic
tech sky130B
magscale 1 2
timestamp 1734110036
<< locali >>
rect 938 1294 1034 1332
rect 996 633 1034 1294
rect 3162 1024 3446 1072
rect 3168 955 3218 1024
rect 2689 926 3218 955
rect 2689 917 3209 926
rect 2154 774 2190 872
rect 2574 774 2616 902
rect 2689 774 2727 917
rect 2790 848 3037 851
rect 3258 848 3294 850
rect 2790 813 3360 848
rect 1186 736 2728 774
rect 1186 734 1802 736
rect 2790 664 2828 813
rect 2946 810 3360 813
rect 2602 626 2828 664
rect 672 82 790 118
rect 754 -598 790 82
rect 2788 44 2912 82
rect 3044 78 3144 80
rect 3258 78 3294 810
rect 3398 646 3446 1024
rect 3044 44 3294 78
rect 2794 -32 2830 44
rect 1618 -70 1914 -36
rect 2516 -70 2830 -32
rect 3108 42 3294 44
rect 3108 -128 3144 42
rect 3258 36 3294 42
rect 2996 -164 3144 -128
rect 3390 -598 3446 646
rect 754 -632 3446 -598
rect 754 -634 3426 -632
<< viali >>
rect 636 82 672 118
<< metal1 >>
rect 592 1346 3436 1432
rect 595 1327 3434 1346
rect 595 888 637 1327
rect 2951 1282 3434 1327
rect 2951 1273 3432 1282
rect 3062 1252 3432 1273
rect 832 1230 2944 1236
rect 686 1186 2944 1230
rect 688 1098 732 1186
rect 832 1178 2944 1186
rect 1204 1135 1258 1136
rect 684 1092 736 1098
rect 1204 1079 1402 1135
rect 1458 1079 1464 1135
rect 1672 1126 2164 1130
rect 2214 1126 2302 1136
rect 2670 1126 2676 1132
rect 1672 1086 2302 1126
rect 2518 1086 2676 1126
rect 684 1034 736 1040
rect 986 1006 992 1058
rect 1044 1006 1050 1058
rect 1204 1016 1258 1079
rect 1672 1076 2164 1086
rect 2214 1056 2302 1086
rect 2670 1080 2676 1086
rect 2728 1080 2734 1132
rect 3354 1122 3432 1252
rect 595 860 834 888
rect 594 846 834 860
rect 594 790 830 846
rect 730 556 830 790
rect 884 730 928 956
rect 1004 812 1032 1006
rect 1830 960 1886 966
rect 1398 941 1450 947
rect 1304 894 1398 936
rect 1726 904 1830 960
rect 1932 924 1938 976
rect 1990 970 1996 976
rect 1990 930 2096 970
rect 1990 924 1996 930
rect 1830 898 1886 904
rect 1398 883 1450 889
rect 1638 812 1678 872
rect 1938 844 1990 924
rect 2240 858 2302 1056
rect 3352 984 3442 1122
rect 2331 976 2389 982
rect 2389 918 2520 976
rect 2331 912 2389 918
rect 3354 874 3432 984
rect 2240 814 2426 858
rect 2936 838 3432 874
rect 1004 784 1680 812
rect 2240 806 2458 814
rect 2936 806 2998 838
rect 3354 836 3432 838
rect 2240 803 3006 806
rect 2240 802 2302 803
rect 2384 782 3006 803
rect 2424 772 3006 782
rect 2894 748 3006 772
rect 3130 784 3182 790
rect 884 686 2720 730
rect 2936 704 2998 748
rect 3130 726 3182 732
rect 870 556 950 560
rect 644 456 950 556
rect 642 410 950 456
rect 644 404 950 410
rect 778 374 830 404
rect 2676 370 2720 686
rect 3135 480 3177 726
rect 2994 418 3292 480
rect 2676 306 2946 370
rect 2676 302 2720 306
rect 612 126 698 140
rect 612 74 628 126
rect 680 74 698 126
rect 612 62 698 74
rect 780 -176 786 -124
rect 838 -128 844 -124
rect 838 -172 1098 -128
rect 838 -176 844 -172
rect 890 -268 942 -172
rect 1408 -176 1886 -132
rect 1670 -306 1676 -301
rect 884 -314 890 -307
rect 876 -352 890 -314
rect 884 -359 890 -352
rect 942 -359 948 -307
rect 1566 -348 1676 -306
rect 1670 -353 1676 -348
rect 1728 -353 1734 -301
rect 2671 -306 2713 235
rect 2844 -68 2850 -12
rect 2906 -68 3006 -12
rect 2627 -348 2713 -306
rect 2460 -438 2466 -386
rect 2518 -438 2524 -386
rect 636 -603 714 -596
rect 636 -665 644 -603
rect 706 -605 714 -603
rect 2671 -605 2713 -348
rect 2799 -481 2805 -423
rect 2863 -481 2941 -423
rect 706 -647 2713 -605
rect 706 -665 714 -647
rect 636 -672 714 -665
<< via1 >>
rect 684 1040 736 1092
rect 1402 1079 1458 1135
rect 992 1006 1044 1058
rect 2676 1080 2728 1132
rect 1398 889 1450 941
rect 1830 904 1886 960
rect 1938 924 1990 976
rect 2331 918 2389 976
rect 3130 732 3182 784
rect 628 118 680 126
rect 628 82 636 118
rect 636 82 672 118
rect 672 82 680 118
rect 628 74 680 82
rect 786 -176 838 -124
rect 890 -359 942 -307
rect 1676 -353 1728 -301
rect 2850 -68 2906 -12
rect 2466 -438 2518 -386
rect 644 -665 706 -603
rect 2805 -481 2863 -423
<< metal2 >>
rect 1005 1409 3319 1447
rect 1005 1332 1043 1409
rect 678 1040 684 1092
rect 736 1040 742 1092
rect 1004 1064 1043 1332
rect 1106 1303 2722 1370
rect 1105 1273 2722 1303
rect 1105 1226 1242 1273
rect 1947 1236 2722 1273
rect 992 1058 1044 1064
rect 688 770 732 1040
rect 992 1000 1044 1006
rect 1105 862 1202 1226
rect 1402 1178 1886 1234
rect 1402 1135 1458 1178
rect 1402 1073 1458 1079
rect 1830 960 1886 1178
rect 1944 1196 2722 1236
rect 1944 982 1984 1196
rect 2682 1138 2722 1196
rect 2676 1132 2728 1138
rect 2676 1074 2728 1080
rect 1938 976 1990 982
rect 1392 889 1398 941
rect 1450 936 1456 941
rect 1450 894 1561 936
rect 1824 904 1830 960
rect 1886 904 1892 960
rect 1938 918 1990 924
rect 2325 918 2331 976
rect 2389 919 2761 976
rect 3281 919 3319 1409
rect 2389 918 3437 919
rect 1450 889 1456 894
rect 1048 810 1202 862
rect 1048 806 1148 810
rect 688 726 834 770
rect 612 130 698 140
rect 612 70 624 130
rect 684 70 698 130
rect 612 62 698 70
rect 790 -118 834 726
rect 1048 68 1104 806
rect 1519 779 1561 894
rect 2703 861 3437 918
rect 3281 859 3319 861
rect 3124 779 3130 784
rect 1519 737 3130 779
rect 3124 732 3130 737
rect 3182 732 3188 784
rect 1048 12 2584 68
rect 2528 -12 2584 12
rect 2850 -12 2906 -6
rect 2528 -68 2850 -12
rect 2850 -74 2906 -68
rect 786 -124 838 -118
rect 786 -182 838 -176
rect 1676 -301 1728 -295
rect 890 -307 942 -301
rect 775 -352 890 -314
rect 775 -539 813 -352
rect 1992 -306 2046 -292
rect 1728 -320 2046 -306
rect 1728 -348 2037 -320
rect 1676 -359 1728 -353
rect 890 -365 942 -359
rect 2466 -386 2518 -380
rect 2466 -444 2518 -438
rect 2805 -423 2863 -417
rect 2473 -539 2511 -444
rect 775 -577 2511 -539
rect 2805 -587 2863 -481
rect 3379 -587 3437 861
rect 636 -603 714 -596
rect 636 -665 644 -603
rect 706 -665 714 -603
rect 2805 -645 3437 -587
rect 636 -672 714 -665
<< via2 >>
rect 624 126 684 130
rect 624 74 628 126
rect 628 74 680 126
rect 680 74 684 126
rect 624 70 684 74
rect 647 -662 703 -606
<< metal3 >>
rect 619 130 689 135
rect 619 70 624 130
rect 684 126 689 130
rect 684 70 1304 126
rect 619 65 1304 70
rect 634 62 1304 65
rect 618 -602 728 -574
rect 618 -666 643 -602
rect 707 -666 728 -602
rect 618 -696 728 -666
<< via3 >>
rect 643 -606 707 -602
rect 643 -662 647 -606
rect 647 -662 703 -606
rect 703 -662 707 -606
rect 643 -666 707 -662
<< metal4 >>
rect 644 -312 1298 -250
rect 644 -601 706 -312
rect 642 -602 708 -601
rect 642 -666 643 -602
rect 707 -666 708 -602
rect 642 -667 708 -666
use N1x1<0.15  N1x1<0.15_0
timestamp 1733686912
transform 1 0 1545 0 1 753
box -53 -53 369 505
use N1x1<0.15  N1x1<0.15_1
timestamp 1733686912
transform 1 0 1123 0 1 753
box -53 -53 369 505
use N1x1<0.15  N1x1<0.15_2
timestamp 1733686912
transform 1 0 1967 0 1 753
box -53 -53 369 505
use N1x1<0.15  N1x1<0.15_3
timestamp 1733686912
transform 1 0 2389 0 1 753
box -53 -53 369 505
use N1x1<1  N1x1<1_0
timestamp 1733623679
transform 1 0 2811 0 1 937
box -53 -53 539 505
use P1x1.5<0.15  P1x1.5<0.15_0
timestamp 1733616804
transform 1 0 701 0 1 753
box -53 -53 369 615
use P1x1<10  P1x1<10_0
timestamp 1733616549
transform 1 0 779 0 1 53
box -53 -53 1979 647
use P1x2<0.15  P1x2<0.15_0
timestamp 1733616004
transform 1 0 2604 0 1 -746
box 154 94 576 862
use P1x2<0.15  P1x2<0.15_1
timestamp 1733616004
transform 1 0 2604 0 1 22
box 154 94 576 862
use P2x7.5<0.15  P2x7.5<0.15_0
timestamp 1733623124
transform 1 0 799 0 1 -599
box -53 -53 953 599
use P2x7.5<0.15  P2x7.5<0.15_1
timestamp 1733623124
transform 1 0 1805 0 1 -599
box -53 -53 953 599
use sky130_fd_pr__cap_mim_m3_1_5Y6EN5  sky130_fd_pr__cap_mim_m3_1_5Y6EN5_0
timestamp 1733670691
transform 1 0 2020 0 1 302
box -880 -734 880 734
<< labels >>
flabel metal1 1918 710 1918 710 0 FreeSans 800 0 0 0 Vm
flabel metal2 s 3410 160 3410 160 0 FreeSans 800 0 0 0 Vout
port 8 nsew
flabel metal1 s 1970 868 1970 868 0 FreeSans 800 0 0 0 I100n
port 11 nsew
flabel metal1 704 466 704 468 0 FreeSans 800 0 0 0 I10n
port 15 nsew
flabel metal1 s 3230 452 3230 452 0 FreeSans 800 0 0 0 Iext
port 19 nsew
flabel locali s 3274 818 3274 818 0 FreeSans 800 0 0 0 Vdd
port 21 nsew
flabel locali s 3336 1048 3336 1048 0 FreeSans 800 0 0 0 Vss
port 23 nsew
<< end >>
