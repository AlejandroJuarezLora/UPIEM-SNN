magic
tech sky130B
magscale 1 2
timestamp 1733620762
<< nwell >>
rect -503 -326 503 326
<< pmos >>
rect -303 -107 -273 107
rect -207 -107 -177 107
rect -111 -107 -81 107
rect -15 -107 15 107
rect 81 -107 111 107
rect 177 -107 207 107
rect 273 -107 303 107
<< pdiff >>
rect -365 95 -303 107
rect -365 -95 -353 95
rect -319 -95 -303 95
rect -365 -107 -303 -95
rect -273 95 -207 107
rect -273 -95 -257 95
rect -223 -95 -207 95
rect -273 -107 -207 -95
rect -177 95 -111 107
rect -177 -95 -161 95
rect -127 -95 -111 95
rect -177 -107 -111 -95
rect -81 95 -15 107
rect -81 -95 -65 95
rect -31 -95 -15 95
rect -81 -107 -15 -95
rect 15 95 81 107
rect 15 -95 31 95
rect 65 -95 81 95
rect 15 -107 81 -95
rect 111 95 177 107
rect 111 -95 127 95
rect 161 -95 177 95
rect 111 -107 177 -95
rect 207 95 273 107
rect 207 -95 223 95
rect 257 -95 273 95
rect 207 -107 273 -95
rect 303 95 365 107
rect 303 -95 319 95
rect 353 -95 365 95
rect 303 -107 365 -95
<< pdiffc >>
rect -353 -95 -319 95
rect -257 -95 -223 95
rect -161 -95 -127 95
rect -65 -95 -31 95
rect 31 -95 65 95
rect 127 -95 161 95
rect 223 -95 257 95
rect 319 -95 353 95
<< nsubdiff >>
rect -467 256 -371 290
rect 371 256 467 290
rect -467 -256 -433 256
rect 433 -256 467 256
rect -467 -290 467 -256
<< nsubdiffcont >>
rect -371 256 371 290
<< poly >>
rect -225 188 -159 204
rect -225 154 -209 188
rect -175 154 -159 188
rect -225 138 -159 154
rect -33 188 33 204
rect -33 154 -17 188
rect 17 154 33 188
rect -33 138 33 154
rect 159 188 225 204
rect 159 154 175 188
rect 209 154 225 188
rect 159 138 225 154
rect -303 107 -273 133
rect -207 107 -177 138
rect -111 107 -81 133
rect -15 107 15 138
rect 81 107 111 133
rect 177 107 207 138
rect 273 107 303 133
rect -303 -138 -273 -107
rect -207 -133 -177 -107
rect -111 -138 -81 -107
rect -15 -133 15 -107
rect 81 -138 111 -107
rect 177 -133 207 -107
rect 273 -138 303 -107
rect -321 -154 -255 -138
rect -321 -188 -305 -154
rect -271 -188 -255 -154
rect -321 -204 -255 -188
rect -129 -154 -63 -138
rect -129 -188 -113 -154
rect -79 -188 -63 -154
rect -129 -204 -63 -188
rect 63 -154 129 -138
rect 63 -188 79 -154
rect 113 -188 129 -154
rect 63 -204 129 -188
rect 255 -154 321 -138
rect 255 -188 271 -154
rect 305 -188 321 -154
rect 255 -204 321 -188
<< polycont >>
rect -209 154 -175 188
rect -17 154 17 188
rect 175 154 209 188
rect -305 -188 -271 -154
rect -113 -188 -79 -154
rect 79 -188 113 -154
rect 271 -188 305 -154
<< locali >>
rect -387 256 -371 290
rect 371 256 387 290
rect -225 154 -209 188
rect -175 154 -159 188
rect -33 154 -17 188
rect 17 154 33 188
rect 159 154 175 188
rect 209 154 225 188
rect -353 95 -319 111
rect -353 -111 -319 -95
rect -257 95 -223 111
rect -257 -111 -223 -95
rect -161 95 -127 111
rect -161 -111 -127 -95
rect -65 95 -31 111
rect -65 -111 -31 -95
rect 31 95 65 111
rect 31 -111 65 -95
rect 127 95 161 111
rect 127 -111 161 -95
rect 223 95 257 111
rect 223 -111 257 -95
rect 319 95 353 111
rect 319 -111 353 -95
rect -321 -188 -305 -154
rect -271 -188 -255 -154
rect -129 -188 -113 -154
rect -79 -188 -63 -154
rect 63 -188 79 -154
rect 113 -188 129 -154
rect 255 -188 271 -154
rect 305 -188 321 -154
<< viali >>
rect -209 154 -175 188
rect -17 154 17 188
rect 175 154 209 188
rect -353 -95 -319 95
rect -257 -57 -223 57
rect -161 -95 -127 95
rect -65 -57 -31 57
rect 31 -95 65 95
rect 127 -57 161 57
rect 223 -95 257 95
rect 319 -57 353 57
rect -305 -188 -271 -154
rect -113 -188 -79 -154
rect 79 -188 113 -154
rect 271 -188 305 -154
<< metal1 >>
rect -221 192 -163 194
rect -29 192 29 194
rect 163 192 221 194
rect -224 188 226 192
rect -224 154 -209 188
rect -175 154 -17 188
rect 17 154 175 188
rect 209 154 226 188
rect -224 142 226 154
rect -359 95 -313 107
rect -359 -95 -353 95
rect -319 -95 -313 95
rect -167 95 -121 107
rect -263 57 -217 69
rect -263 -57 -257 57
rect -223 -57 -217 57
rect -263 -69 -217 -57
rect -359 -107 -313 -95
rect -167 -95 -161 95
rect -127 -95 -121 95
rect 25 95 71 107
rect -71 57 -25 69
rect -71 -57 -65 57
rect -31 -57 -25 57
rect -71 -69 -25 -57
rect -167 -107 -121 -95
rect 25 -95 31 95
rect 65 -95 71 95
rect 217 95 263 107
rect 121 57 167 69
rect 121 -57 127 57
rect 161 -57 167 57
rect 121 -69 167 -57
rect 25 -107 71 -95
rect 217 -95 223 95
rect 257 -95 263 95
rect 313 57 359 69
rect 313 -57 319 57
rect 353 -57 359 57
rect 313 -69 359 -57
rect 217 -107 263 -95
rect -317 -154 -259 -148
rect -317 -176 -305 -154
rect -322 -188 -305 -176
rect -271 -176 -259 -154
rect -125 -154 -67 -148
rect -125 -176 -113 -154
rect -271 -188 -113 -176
rect -79 -176 -67 -154
rect 67 -154 125 -148
rect 67 -176 79 -154
rect -79 -188 79 -176
rect 113 -176 125 -154
rect 259 -154 317 -148
rect 259 -176 271 -154
rect 113 -188 271 -176
rect 305 -188 317 -154
rect -322 -194 317 -188
rect -322 -228 316 -194
<< properties >>
string FIXED_BBOX -450 -273 450 273
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.07 l 0.15 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 60 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
