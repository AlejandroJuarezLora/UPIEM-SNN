** sch_path: /home/ashley/Desktop/Modelo_Neronal_1/NeuronaFinal.sch
.subckt NeuronaFinal Vout I100n Vdd Vss Iext I10n
*.PININFO Vout:B I100n:B Vdd:B Vss:B Iext:B I10n:B
XM1 I10n I10n Vm Vdd sky130_fd_pr__pfet_01v8 L=10 W=1 nf=1 m=1
XM2 Vm net1 I10n Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=1.5 nf=1 m=1
XM3 net1 net1 Vm Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=7.5 nf=1 m=2
XM4 net1 I10n Vss Vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM5 I100n I10n Vss Vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM6 Vout I100n Vdd Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM7 Vout I100n Vss Vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XM8 net2 net2 Iext Vss sky130_fd_pr__nfet_01v8 L=1 W=1 nf=1 m=1
XM9 Vm I10n Iext Vdd sky130_fd_pr__pfet_01v8 L=0.15 W=2 nf=1 m=1
XM10 Vout I10n net2 Vss sky130_fd_pr__nfet_01v8 L=0.15 W=1 nf=1 m=1
XC1 Vm Vss sky130_fd_pr__cap_mim_m3_1 W=22 L=23 m=1
.ends
.end
