magic
tech sky130B
magscale 1 2
timestamp 1733623124
<< nwell >>
rect -503 -326 503 326
<< pmos >>
rect -303 -107 -273 107
rect -207 -107 -177 107
rect -111 -107 -81 107
rect -15 -107 15 107
rect 81 -107 111 107
rect 177 -107 207 107
rect 273 -107 303 107
<< pdiff >>
rect -365 95 -303 107
rect -365 -95 -353 95
rect -319 -95 -303 95
rect -365 -107 -303 -95
rect -273 95 -207 107
rect -273 -95 -257 95
rect -223 -95 -207 95
rect -273 -107 -207 -95
rect -177 95 -111 107
rect -177 -95 -161 95
rect -127 -95 -111 95
rect -177 -107 -111 -95
rect -81 95 -15 107
rect -81 -95 -65 95
rect -31 -95 -15 95
rect -81 -107 -15 -95
rect 15 95 81 107
rect 15 -95 31 95
rect 65 -95 81 95
rect 15 -107 81 -95
rect 111 95 177 107
rect 111 -95 127 95
rect 161 -95 177 95
rect 111 -107 177 -95
rect 207 95 273 107
rect 207 -95 223 95
rect 257 -95 273 95
rect 207 -107 273 -95
rect 303 95 365 107
rect 303 -95 319 95
rect 353 -95 365 95
rect 303 -107 365 -95
<< pdiffc >>
rect -353 -95 -319 95
rect -257 -95 -223 95
rect -161 -95 -127 95
rect -65 -95 -31 95
rect 31 -95 65 95
rect 127 -95 161 95
rect 223 -95 257 95
rect 319 -95 353 95
<< nsubdiff >>
rect -467 256 -371 290
rect 371 256 467 290
rect -467 -256 -433 256
rect 433 -256 467 256
rect -467 -290 467 -256
<< nsubdiffcont >>
rect -371 256 371 290
<< poly >>
rect -225 188 -159 204
rect -225 154 -209 188
rect -175 154 -159 188
rect -225 138 -159 154
rect -33 188 33 204
rect -33 154 -17 188
rect 17 154 33 188
rect -33 138 33 154
rect 159 188 225 204
rect 159 154 175 188
rect 209 154 225 188
rect 159 138 225 154
rect -303 107 -273 133
rect -207 107 -177 138
rect -111 107 -81 133
rect -15 107 15 138
rect 81 107 111 133
rect 177 107 207 138
rect 273 107 303 133
rect -303 -138 -273 -107
rect -207 -133 -177 -107
rect -111 -138 -81 -107
rect -15 -133 15 -107
rect 81 -138 111 -107
rect 177 -133 207 -107
rect 273 -138 303 -107
rect -321 -154 -255 -138
rect -321 -188 -305 -154
rect -271 -188 -255 -154
rect -321 -204 -255 -188
rect -129 -154 -63 -138
rect -129 -188 -113 -154
rect -79 -188 -63 -154
rect -129 -204 -63 -188
rect 63 -154 129 -138
rect 63 -188 79 -154
rect 113 -188 129 -154
rect 63 -204 129 -188
rect 255 -154 321 -138
rect 255 -188 271 -154
rect 305 -188 321 -154
rect 255 -204 321 -188
<< polycont >>
rect -209 154 -175 188
rect -17 154 17 188
rect 175 154 209 188
rect -305 -188 -271 -154
rect -113 -188 -79 -154
rect 79 -188 113 -154
rect 271 -188 305 -154
<< locali >>
rect -387 256 -371 290
rect 371 256 387 290
rect -225 154 -209 188
rect -175 154 -159 188
rect -33 154 -17 188
rect 17 154 33 188
rect 159 154 175 188
rect 209 154 225 188
rect -353 95 -319 111
rect -353 -111 -319 -95
rect -257 95 -223 111
rect -257 -111 -223 -95
rect -161 95 -127 111
rect -161 -111 -127 -95
rect -65 95 -31 111
rect -65 -111 -31 -95
rect 31 95 65 111
rect 31 -111 65 -95
rect 127 95 161 111
rect 127 -111 161 -95
rect 223 95 257 111
rect 223 -111 257 -95
rect 319 95 353 111
rect 319 -111 353 -95
rect -321 -188 -305 -154
rect -271 -188 -255 -154
rect -129 -188 -113 -154
rect -79 -188 -63 -154
rect 63 -188 79 -154
rect 113 -188 129 -154
rect 255 -188 271 -154
rect 305 -188 321 -154
<< viali >>
rect -209 154 -175 188
rect -17 154 17 188
rect 175 154 209 188
rect -353 -95 -319 95
rect -257 -48 -223 48
rect -161 -95 -127 95
rect -65 -48 -31 48
rect 31 -95 65 95
rect 127 -48 161 48
rect 223 -95 257 95
rect 319 -48 353 48
rect -305 -188 -271 -154
rect -113 -188 -79 -154
rect 79 -188 113 -154
rect 271 -188 305 -154
<< metal1 >>
rect -224 188 226 198
rect -224 184 -209 188
rect -472 154 -209 184
rect -175 154 -17 188
rect 17 154 175 188
rect 209 154 226 188
rect -472 152 226 154
rect -472 -168 -440 152
rect -224 146 226 152
rect -359 95 -313 107
rect -359 -95 -353 95
rect -319 -92 -313 95
rect -167 95 -121 107
rect -263 48 -217 60
rect -263 25 -257 48
rect -223 31 -217 48
rect -223 25 -210 31
rect -263 -27 -262 25
rect -263 -48 -257 -27
rect -223 -33 -210 -27
rect -223 -48 -217 -33
rect -263 -60 -217 -48
rect -167 -92 -161 95
rect -319 -95 -161 -92
rect -127 -92 -121 95
rect 25 95 71 107
rect -71 48 -25 60
rect -71 31 -65 48
rect -74 25 -65 31
rect -31 31 -25 48
rect -31 25 -22 31
rect -74 -33 -65 -27
rect -71 -48 -65 -33
rect -31 -33 -22 -27
rect -31 -48 -25 -33
rect -71 -60 -25 -48
rect 25 -92 31 95
rect -127 -95 31 -92
rect 65 -92 71 95
rect 217 95 263 107
rect 121 48 167 60
rect 121 31 127 48
rect 118 25 127 31
rect 161 31 167 48
rect 161 25 170 31
rect 118 -33 127 -27
rect 121 -48 127 -33
rect 161 -33 170 -27
rect 161 -48 167 -33
rect 121 -60 167 -48
rect 217 -92 223 95
rect 65 -95 223 -92
rect 257 -90 263 95
rect 313 48 359 60
rect 313 25 319 48
rect 353 25 359 48
rect 306 -27 312 25
rect 364 20 370 25
rect 364 -22 414 20
rect 364 -27 370 -22
rect 313 -48 319 -27
rect 353 -48 359 -27
rect 313 -60 359 -48
rect 257 -95 264 -90
rect -359 -107 264 -95
rect -358 -120 264 -107
rect -317 -154 -259 -148
rect -317 -156 -305 -154
rect -322 -168 -305 -156
rect -472 -188 -305 -168
rect -271 -156 -259 -154
rect -125 -154 -67 -148
rect -125 -156 -113 -154
rect -271 -188 -113 -156
rect -79 -156 -67 -154
rect 67 -154 125 -148
rect 67 -156 79 -154
rect -79 -188 79 -156
rect 113 -156 125 -154
rect 259 -154 317 -148
rect 259 -156 271 -154
rect 113 -188 271 -156
rect 305 -156 317 -154
rect 305 -188 322 -156
rect -472 -200 322 -188
rect -322 -204 322 -200
<< via1 >>
rect -262 -27 -257 25
rect -257 -27 -223 25
rect -223 -27 -210 25
rect -74 -27 -65 25
rect -65 -27 -31 25
rect -31 -27 -22 25
rect 118 -27 127 25
rect 127 -27 161 25
rect 161 -27 170 25
rect 312 -27 319 25
rect 319 -27 353 25
rect 353 -27 364 25
<< metal2 >>
rect 312 25 364 31
rect -268 -27 -262 25
rect -210 20 -204 25
rect -80 20 -74 25
rect -210 -22 -74 20
rect -210 -27 -204 -22
rect -80 -27 -74 -22
rect -22 20 -16 25
rect 112 20 118 25
rect -22 -22 118 20
rect -22 -27 -16 -22
rect 112 -27 118 -22
rect 170 20 176 25
rect 170 -22 312 20
rect 170 -27 176 -22
rect 312 -33 364 -27
<< labels >>
flabel metal1 s 0 170 0 170 0 FreeSans 320 0 0 0 G
port 0 nsew
flabel metal1 s -338 -2 -338 -2 0 FreeSans 320 0 0 0 D
port 1 nsew
flabel metal1 s 388 0 388 0 0 FreeSans 320 0 0 0 S
port 2 nsew
flabel locali s -18 274 -18 274 0 FreeSans 320 0 0 0 B
port 4 nsew
<< properties >>
string FIXED_BBOX -450 -273 450 273
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.07 l 0.15 m 1 nf 7 diffcov 100 polycov 100 guard 1 glc 0 grc 0 gtc 1 gbc 0 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 0 viasrc 50 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
