magic
tech sky130B
magscale 1 2
timestamp 1733686912
use sky130_fd_pr__nfet_01v8_RZ9R45  sky130_fd_pr__nfet_01v8_RZ9R45_0
timestamp 1733686912
transform 1 0 158 0 1 226
box -211 -279 211 279
<< end >>
